module channel_module(input clk, rst, SW1, SW2, add, input[3:0] address, data, input valid, output ack, output[3:0] data_out, output data_out_valid, output[1:0] channel, output channel_valid);
    
endmodule